// Verilog netlist created by TD v4.6.18154
// Wed Apr 29 19:53:00 2020

`timescale 1ns / 1ps
module sysmem_mh  // al_ip/mem_mh/mem_mh.v(14)
  (
  addra,
  cea,
  clka,
  dia,
  wea,
  doa
  );

  input [9:0] addra;  // al_ip/mem_mh/mem_mh.v(19)
  input cea;  // al_ip/mem_mh/mem_mh.v(21)
  input clka;  // al_ip/mem_mh/mem_mh.v(22)
  input [7:0] dia;  // al_ip/mem_mh/mem_mh.v(18)
  input wea;  // al_ip/mem_mh/mem_mh.v(20)
  output [7:0] doa;  // al_ip/mem_mh/mem_mh.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h413E93830007F1B78993830001228272E5F707F1B7E7F4C1B7A3000120010000),
    .INIT_01(256'h72C4F98323038444BA03832344252323232282220107C48507E417C419232279),
    .INIT_02(256'h2201C00113800006823285E3830323C429F707B6838303C4C405232323232282),
    .INIT_03(256'h068262013E8304BD833E8304F79183232393B72393B72393B72393B7A3800682),
    .INIT_04(256'h833E938411133E93833E93441DF7C1833E9344811323832323227941B2213100),
    .INIT_05(256'h83007907BA0383005DF7444DF7A1833E9344F9F7E183F4BA8303BD83048D3E93),
    .INIT_06(256'h525000E7F7E10323843123A3F4E7F4000D2350E1B7A323223945B2F784C4F485),
    .INIT_07(256'h2069786F79656D000D656E637700726C6531720A3832456F616E6E7541433320),
    .INIT_08(256'h000000000000000000000000000000000000000000000000000000002E552047),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_1024x8_sub_000000_000 (
    .addra({addra,3'b111}),
    .cea(cea),
    .clka(clka),
    .dia({open_n68,dia}),
    .wea(wea),
    .doa({open_n83,doa}));

endmodule 

